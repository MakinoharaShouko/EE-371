module new_object (old_queue, clk, new_queue);
	input logic clk;
	input object[] old_queue;
	output object[] new_queue;
endmodule
