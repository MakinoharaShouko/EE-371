module DE1_SoC (CLOCK_50);
	input logic CLOCK_50;
	
	object o [$] = {};
endmodule
